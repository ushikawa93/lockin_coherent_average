
module clocks (
	clk_clk,
	clk_ca_clk,
	clk_calc_finales_clk,
	clk_lockin_clasico_clk,
	clk_ma_clk,
	reset_reset_n);	

	input		clk_clk;
	output		clk_ca_clk;
	output		clk_calc_finales_clk;
	output		clk_lockin_clasico_clk;
	output		clk_ma_clk;
	input		reset_reset_n;
endmodule
