// clocks.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module clocks (
		input  wire  clk_clk,           //           clk.clk
		output wire  clk_lento_clk,     //     clk_lento.clk
		output wire  clk_mas_lento_clk, // clk_mas_lento.clk
		output wire  clk_rapido_clk,    //    clk_rapido.clk
		input  wire  reset_reset_n      //         reset.reset_n
	);

	clocks_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (clk_rapido_clk),    // outclk0.clk
		.outclk_1 (clk_lento_clk),     // outclk1.clk
		.outclk_2 (clk_mas_lento_clk), // outclk2.clk
		.locked   ()                   // (terminated)
	);

endmodule
