// clocks.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module clocks (
		input  wire  clk_clk,                //                clk.clk
		output wire  clk_ca_clk,             //             clk_ca.clk
		output wire  clk_calc_finales_clk,   //   clk_calc_finales.clk
		output wire  clk_lockin_clasico_clk, // clk_lockin_clasico.clk
		output wire  clk_ma_clk,             //             clk_ma.clk
		input  wire  reset_reset_n           //              reset.reset_n
	);

	clocks_pll_0 pll_0 (
		.refclk   (clk_clk),                //  refclk.clk
		.rst      (~reset_reset_n),         //   reset.reset
		.outclk_0 (clk_lockin_clasico_clk), // outclk0.clk
		.outclk_1 (clk_ca_clk),             // outclk1.clk
		.outclk_2 (clk_ma_clk),             // outclk2.clk
		.outclk_3 (clk_calc_finales_clk),   // outclk3.clk
		.locked   ()                        // (terminated)
	);

endmodule
